/*package i2c_vip_package;

`include "uvm_macros.svh"

import uvm_pkg::*;



//`include "apb_seq_item.sv"
`include "i2c_slave_tx_item.sv"


`include "apb_config_obj.sv"
`include "i2c_slave_config.sv"
`include "i2c_env_config.sv"

//`include "apb_sequencer.sv"
`include "apb_driver.sv"
`include "apb_monitor.sv"
`include "apb_agent.sv"
`include "apb_sequence.sv"
`include "wr_rd_seq.sv"
`include "apb_seq_item.sv"
//`include "apb_reset_seq.sv"


`include "i2c_slave_sequencer.sv"
`include "i2c_slave_driver.sv"
`include "i2c_slave_monitor.sv"
`include "i2c_slave_agent.sv"

`include "i2c_vip_scoreboard.sv"
`include "i2c_vip_env.sv"

//`include "i2c_seqs.sv"




`include "i2c_vip_test.sv"
//`include "i2c_apb_vip_reset_test.sv"
`include "i2c_apb_vip_wr_rd_test.sv"


endpackage */
